`include "define.v"

module InitMap (
    input reset,
    output reg [`tile_col_num * `tile_row_num - 1:0] tilemap_dots,
    output reg [`tile_col_num * `tile_row_num - 1:0] tilemap_big_dots
);

    // wire [`tile_col_num * `tile_row_num - 1:0] init_dots;
    // wire [`tile_col_num * `tile_row_num - 1:0] init_big_dots;

    // integer i;
    // reg [`tile_col_num - 1:0] temp [0: `tile_row_num - 1];

    // initial begin
        // $readmemb("./maps/walls.txt", temp);
        // for (i = 0; i < `tile_row_num; i = i + 1) begin
        //     init_walls[i * `tile_col_num +: `tile_col_num] = temp[i];
        // end
        // $readmemb("./maps/dots.txt", temp);
        // for (i = 0; i < `tile_row_num; i = i + 1) begin
        //     init_dots[i * `tile_col_num +: `tile_col_num] = temp[i];
        // end
        // $readmemb("./maps/big_dots.txt", temp);
        // for (i = 0; i < `tile_row_num; i = i + 1) begin
        //     init_big_dots[i * `tile_col_num +: `tile_col_num] = temp[i];
        // end
    // end

    always @(negedge reset) begin
        tilemap_dots <=     768'b000000000000000000000000000000000111111110111100001111111111111001000001000001000010000010000010010000010000010000100000100000100111111111111111111111111111111001000001001000000000010010000010010000010010000000000100100000100111111100111110011111001111111000000001000000100100000010000000000000010011111111111100100000000000000100100000000001001000000000000001111011111111011110000000000000010010000000000100100000000000000100111111111111001000000000000001001000000000010010000000011111111111111001111111111111100100000100000010010000001000001001111001111111111111111110011110000010010010000000000100100100000000100100100000000001001001000001111111001111100111110011111110010000000000001001000000000000100111111111111111111111111111111000000000000000000000000000000000;
        tilemap_big_dots <= 768'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end

endmodule